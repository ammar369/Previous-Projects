module byte_gen
(
input start,
input [7:0] data_i,		//value in register i
input [7:0] data_j,		//value in register j
input [4:0] data_k,		//value of 5 bit counter register k
input loop_signal,		//for detecting k overflow
input [7:0] ram_data,	//data output by ram and read in

output logic [7:0] data_to_ram,		//data to be sent to ram
output logic [7:0] address_to_ram,	//address to be read from/ or written to
output logic ram_wren,				//tells if we are writing or reading from ram

output logic [7:0] init_count_k,	//initialized value of counter_reg k
output logic start_count_k,			//enables counting of k
output logic pause_k,				//if high, it pauses k, if low, unpauses k

output logic [7:0] reg_in_i,		//input to reg i
output logic reg_enable_i,			//writing to reg i

output logic [7:0] reg_in_j,		//input to reg j
output logic reg_enable_j,			//writing to reg j

output logic [7:0] gen_byte,		//this holds output that we need to get/ f

output logic finish
);

localparam idle 		= 4'b0000;
localparam incrmnt_i 	= 4'b0001;
localparam get_var 		= 4'b0011;
localparam j_read_Sj 	= 4'b0010;
localparam write_Si		= 4'b0110;
localparam write_Sj 	= 4'b0100;
localparam byte_gen		= 4'b0101;
localparam incrmnt_k 	= 4'b0111;
localparam finished 	= 4'b1111;

logic [3:0] state = idle;
logic [3:0] next_state;


logic [7:0] temp_Si;
logic [7:0] temp_j;
logic [7:0] temp_Sj;
logic [7:0] temp_addr;
logic [7:0] temp_f;

always @(posedge clk or posedge reset)
begin
	if (reset) state <= idle;
	else state <= next_state;	
end

always @(*)
begin
	case(state)
	idle:		begin	data_to_ram = 0;
						address_to_ram = 0;
						ram_wren = 0;
						init_count_k = 0;
						start_count_k = 0;
						pause_k = 0;
						reg_in_i = 0;
						reg_enable_i = 0;
						reg_in_j = 0;
						reg_enable_j = 0;
						next_state <= start ? get_var : idle;		//if start is high, we start operation
				end
	incrmnt_i:	begin	pause_k = 1'b1;								//pauses value of k so that we can compute for that value
						if (loop_signal) next_state <= finished;	//loop signal tells if i overflows (reaches 256) and it then stops the loop
						temp_i <= data_i + 1'b1;	//value of i is incremented and passed to temp_i
						reg_in_i = temp_i;			//temp_i overwrites old value of i
						reg_enable_i = 1'b1;		//writing to reg_i enabled
						address_to_ram <= temp_i;	//we get value at incremented i S[i+1]
						next_state <= get_var;
				end
	get_var:	begin	temp_Si = ram_data;			//data from ram is stored in a temp variable
						temp_j = data_j + ram_data	//we take in old value of j, and S[i](in ram data) to get new value of j
						next_state <= j_read_Sj;
				end
	j_read_Sj:	begin	reg_in = temp_j;			//we update value of j stored in register
						reg_enable = 1'b1;			//we write to register with new j
						address_to_ram <= temp_j;	//we read S[j]
						next_state <= write_Si;
				end
	write_Si:	begin	temp_Sj = ram_data;			//S[j] is stored in variable
						data_to_ram = temp_Sj;		//S[j] is data to be written in ram
						address_to_ram = data_i;	//it is to be written at address of i, so S[i] = S[j]
						ram_wren = 1'b1;			//we start writing
						next_state <= write_Sj;
				end
	write_Sj:	begin	data_to_ram = temp_Si;		//we take value of S[i] and send that to be written to ram
						address_to_ram = data_j;	//we write the data at address S[j]
						ram_wren = 1'b1;			
						temp_addr = temp_Si + temp_Sj;
						address_to_ram = temp_addr;
						next_state <= byte_gen;
				end
	byte_gen:	begin	temp_f = ram_data;			//we get f from the address computed
						gen_byte = temp_f;			//we update output to give the generated byte
						next_state <= incrmnt_k;
				end
	incrmnt_k:	begin	start_count_k = 1'b1;		//we start k counter (if for first time, k=0)
						pause_k = 1'b0;				//we unpause k counter for subsequent times
						next_state <= incrmnt_i;	//we restart loop
				end
	finished:	begin	finish = 1;					//when loop computes 256 times, we finish execution
						next_state <= idle;			//then we again go to idle state to wait for next start input
				end
	default:	next_state <= idle;
	endcase
end

endmodule